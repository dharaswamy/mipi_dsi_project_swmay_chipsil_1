
//----------------------------------------------------------
//
//----------------------------------------------------------


//---------------------------------------------------------------------------------------------------------
class pxl_config_agent extends uvm_object;
  
//factory registration.
  `uvm_object_utils(pxl_config_agent)
  
  uvm_active_passive_enum is_active = UVM_ACTIVE ;
  
  function new(string name = "pxl_config_agent");
    super.new(name);
    `uvm_info("TRACE",$sformatf("%m"),UVM_HIGH)
  endfunction:new
  
endclass:pxl_config_agent

//----------------------------------------------------------
//
//----------------------------------------------------------


//----------------------------------------------------------
//
//----------------------------------------------------------


//=========================================================================================================