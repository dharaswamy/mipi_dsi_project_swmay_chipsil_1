
//-------------------------------------------------------------------
// Class Name : pxl_monitor
// Type       : uvm_component type
//-------------------------------------------------------------------


//-------------------------------------------------------------------------------------------------------------------

class pxl_monitor extends uvm_monitor;
  
//---------------------------------------------------------------
// Factory registration
// This class is uvm component class so use component_utils_begin
//--------------------------------------------------------------
  `uvm_component_utils(pxl_monitor)
  
//---------------------------------------------------------
// Port type : analysis port
// Usage / purpose  : Sending the transactions to the scoreboard and functional coverage
//---------------------------------------------------------
  uvm_analysis_port#(pxl_sequ_item) 

//---------------------------------------------------------
//
//---------------------------------------------------------


//---------------------------------------------------------
//
//---------------------------------------------------------


//---------------------------------------------------------
//
//---------------------------------------------------------


endclass:pxl_monitor

//===================================================================================================================